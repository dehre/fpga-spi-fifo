package custom_types is

    -- Enumerated type for decimal digits (0-9)
    type t_decimal_digit is (ZERO, ONE, TWO, THREE, FOUR, FIVE, SIX, SEVEN, EIGHT, NINE);

end package;
